
module debugger (
	probe);	

	input	[31:0]	probe;
endmodule
