
module probes (
	source,
	probe);	

	output	[0:0]	source;
	input	[31:0]	probe;
endmodule
